package ca12_dat_130 is

constant ca12_type130:integer:=1;
constant ca12_inve130:integer:=2;
signal ca12_ord130:real_vector(1 to 3):=(4.0, 3.0, 0.0);
signal ca12_fak130:real_vector(1 to 4):=(0.975294676147E-01, 0.220185632619, 0.00000000000, 25.6028993526);
constant ca12_anz130:integer:=       20;
signal ca12_data130:real_vector(1 to 20):=
(
  0.712086240885    ,
  0.186297166892    ,
 -0.208887154143E-01,
  0.531007092724E-02,
 -0.181480706895E-02,
  0.128558883926    ,
 -0.939139994662E-02,
  0.372136915760E-02,
 -0.259077537559E-02,
  0.104687708202E-02,
 -0.293936530550E-02,
  0.667614364241E-03,
 -0.506853279164E-03,
  0.113773216487E-02,
 -0.947577210652E-03,
  0.196412408079E-03,
  0.637444737511E-04,
 -0.129103797161E-03,
 -0.532315735795E-03,
  0.644951605279E-03
);

end;
