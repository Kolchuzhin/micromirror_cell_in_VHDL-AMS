package ca13_dat_130 is

constant ca13_type130:integer:=1;
constant ca13_inve130:integer:=2;
signal ca13_ord130:real_vector(1 to 3):=(4.0, 3.0, 0.0);
signal ca13_fak130:real_vector(1 to 4):=(0.975294676147E-01, 0.220185632619, 0.00000000000, 25.6030000457);
constant ca13_anz130:integer:=       20;
signal ca13_data130:real_vector(1 to 20):=
(
  0.712094286463    ,
 -0.186347802870    ,
 -0.209412180795E-01,
 -0.523557199207E-02,
 -0.178345484280E-02,
  0.128565735753    ,
  0.931339715905E-02,
  0.363612109234E-02,
  0.264112674223E-02,
  0.111307000174E-02,
 -0.294786738552E-02,
 -0.533796708169E-03,
 -0.463952089322E-03,
 -0.131455480646E-02,
 -0.989450152969E-03,
  0.190516958085E-03,
  0.124293432457E-04,
 -0.498349836548E-04,
  0.494604396684E-03,
  0.599958313911E-03
);

end;
