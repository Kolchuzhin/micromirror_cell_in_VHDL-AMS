package s_dat_135 is

constant s_type135:integer:=1;
constant s_inve135:integer:=1;
signal s_ord135:real_vector(1 to 3):=( 6.0, 4.0, 2.0);
signal s_fak135:real_vector(1 to 4):=( 0.985831178093E-01, 0.214896594093, 4.92915589046, 18455.91307);
constant s_anz135:integer:=       105;
signal s_data135:real_vector(1 to 105):=
(
 -0.380462328309E-11,
  0.217133727115E-12,
  0.477269987897    ,
 -0.826024419409E-12,
  0.148695432725E-09,
  0.627133609178E-12,
 -0.172249760625E-09,
  0.703729843662E-14,
 -0.912518157304E-10,
 -0.128631124369E-12,
  0.529133596581E-09,
  0.340831468502E-12,
 -0.434350889708E-09,
 -0.220774222723E-12,
  0.516065208620    ,
 -0.182053570831E-11,
 -0.118904595638E-08,
  0.698466661345E-11,
  0.338750270261E-08,
 -0.531987677792E-11,
 -0.330044812007E-08,
 -0.846830662014E-14,
  0.912589476182E-10,
  0.150556580628E-12,
 -0.529160390626E-09,
 -0.395415686133E-12,
  0.434371027913E-09,
  0.254970913913E-12,
 -0.587993396505E-10,
  0.163107328614E-11,
 -0.105484446381E-08,
 -0.627031540115E-11,
  0.307369937992E-08,
  0.477947544796E-11,
 -0.116531481782E-08,
  0.179176936707E-15,
 -0.144754500760E-10,
 -0.314523523583E-14,
  0.203752572084E-09,
  0.793546415820E-14,
 -0.189940194776E-09,
 -0.498992950459E-14,
 -0.293910389349E-10,
 -0.746235378567E-23,
  0.866197505189E-10,
  0.208035814297E-22,
 -0.665457030012E-10,
 -0.128033527996E-22,
  0.922414811689E-11,
 -0.895884802457E-15,
  0.231259325235E-09,
  0.157261783745E-13,
 -0.146606319931E-08,
 -0.396773266580E-13,
  0.123912979062E-08,
  0.249496513426E-13,
  0.119169846151E-10,
  0.619056888255E-23,
  0.124994753643E-10,
 -0.148198281620E-22,
 -0.981768325965E-10,
  0.784802677662E-23,
  0.737751906659E-10,
  0.716707869137E-15,
 -0.216783893369E-09,
 -0.125809432015E-13,
  0.126231079439E-08,
  0.317418626682E-13,
 -0.104918976477E-08,
 -0.199597219479E-13,
  0.666480376456E-02,
 -0.213631186640E-12,
 -0.113633752522E-10,
  0.803411496331E-12,
 -0.144999700034E-09,
 -0.606899569818E-12,
  0.161665008295E-09,
 -0.189178829934E-14,
  0.170703658697E-09,
  0.322788514369E-13,
 -0.752822985110E-09,
 -0.799608870022E-13,
  0.579094210710E-09,
  0.497468720851E-13,
 -0.661965555697E-10,
  0.178983745133E-11,
  0.991354764861E-09,
 -0.680335546375E-11,
 -0.268453764737E-08,
  0.516054891875E-11,
  0.202646318583E-08,
  0.257670397685E-14,
 -0.170711122996E-09,
 -0.400978138646E-13,
  0.752850963234E-09,
  0.963143724992E-13,
 -0.579115225064E-09,
 -0.588587644605E-13,
  0.473064745010E-10,
 -0.160275186343E-11,
 -0.458177827975E-09,
  0.610677897394E-11,
  0.186371332836E-08,
 -0.463650995299E-11,
 -0.166566309091E-08
);
end;
