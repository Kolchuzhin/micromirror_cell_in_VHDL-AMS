package initial is

constant mm_1:real:=  0.287950035810E-08;
constant dm_1:real:=  0.702143607267E-04;
constant mm_2:real:=  0.659733846875E-08;
constant dm_2:real:=  0.240906751644E-03;
constant mm_3:real:=  0.263744816095E-08;
constant dm_3:real:=  0.397046131356E-03;
constant fi1_1:real:= -0.997749461172    ;
constant fi1_2:real:=  0.999999999998    ;
constant fi1_3:real:= -0.714154416552    ;
constant fi2_1:real:=  0.215667880024E-10;
constant fi2_2:real:=  0.996525353204    ;
constant fi2_3:real:= -0.705805491469    ;
constant fi3_1:real:=  0.997749461215    ;
constant fi3_2:real:=  0.999999999883    ;
constant fi3_3:real:= -0.714154416561    ;
constant el1_1:real:=  0.141920120004E-11;
constant el1_2:real:= -0.709831408332E-01;
constant el1_3:real:= -0.317009944282E-02;
constant el2_1:real:=  -60732.3144099    ;
constant el2_2:real:=   103560.713601    ;
constant el2_3:real:=   4625.29581182    ;                        
end;
