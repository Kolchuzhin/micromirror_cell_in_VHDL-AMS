package ca23_dat_130 is

constant ca23_type130:integer:=1;
constant ca23_inve130:integer:=2;
signal ca23_ord130:real_vector(1 to 3):=(4.0, 3.0, 0.0);
signal ca23_fak130:real_vector(1 to 4):=(0.975294676147E-01, 0.220185632619, 0.00000000000, 4353.18490300);
constant ca23_anz130:integer:=       20;
signal ca23_data130:real_vector(1 to 20):=
(
  0.546111390319    ,
  0.295871790946E-03,
  0.879069075222E-02,
 -0.293891270388E-03,
 -0.641224996279E-03,
 -0.263461122282    ,
 -0.718573965052E-03,
 -0.864593553516E-03,
  0.173269568371E-02,
 -0.516914738996E-02,
  0.125610539761    ,
 -0.128446242254E-02,
  0.499953901998E-02,
  0.127235001362E-02,
 -0.131318972091E-02,
 -0.444623172071E-01,
  0.163315957039E-02,
 -0.909045625811E-02,
 -0.260866762118E-02,
  0.702268147666E-02
);

end;
