package ca12_dat_135 is

constant ca12_type135:integer:=1;
constant ca12_inve135:integer:=2;
signal ca12_ord135:real_vector(1 to 3):=( 6.0, 4.0, 2.0);
signal ca12_fak135:real_vector(1 to 4):=( 0.985831178093E-01, 0.214896594093, 4.92915589046, 25.8957269075);
constant ca12_anz135:integer:=       105;
signal ca12_data135:real_vector(1 to 105):=
(
  0.712855361891    ,
 -0.181346587868    ,
 -0.198015186198E-01,
 -0.415927375416E-02,
 -0.153573430027E-02,
 -0.510237922820E-03,
 -0.764100630283E-04,
  0.131880723107    ,
  0.964664849709E-02,
  0.397724201981E-02,
  0.162623410076E-02,
 -0.132542281553E-03,
  0.485582696654E-03,
  0.737744039164E-03,
 -0.307644645158E-02,
 -0.907572318294E-03,
 -0.875589375186E-03,
 -0.202386662848E-03,
  0.233665775380E-03,
 -0.466458263355E-03,
 -0.467484331887E-03,
  0.217954553170E-03,
  0.776231117698E-04,
 -0.997658717706E-04,
 -0.938691903505E-04,
  0.556966054463E-03,
  0.549523243109E-03,
  0.548273297425E-04,
 -0.231063812390E-04,
 -0.525968371687E-04,
 -0.707438293504E-04,
  0.292791303765E-03,
  0.322200008401E-03,
 -0.505699831991E-03,
 -0.530082698612E-03,
  0.421071642029E-03,
  0.152590653211E-03,
  0.295736663012E-04,
  0.117431331453E-04,
  0.766868969508E-05,
  0.527054350921E-05,
  0.166617512612E-05,
  0.445482327591E-04,
  0.358221111798E-04,
  0.432190474514E-04,
 -0.469647211899E-04,
 -0.145540033912E-03,
  0.395419458803E-04,
  0.120682124213E-03,
 -0.268652436678E-04,
 -0.370734016171E-04,
 -0.656911565201E-04,
  0.126956731874E-03,
  0.228073073747E-03,
 -0.129165674348E-03,
 -0.184322337900E-03,
  0.877033943448E-05,
 -0.851429208706E-06,
 -0.476767509670E-04,
  0.366154716279E-04,
  0.225448526368E-03,
 -0.446961499914E-05,
 -0.186547357241E-03,
 -0.299619802769E-05,
  0.262681936434E-04,
  0.532746472007E-04,
 -0.175669246799E-03,
 -0.219657099111E-03,
  0.167451751873E-03,
  0.152887349480E-03,
 -0.219837737744E-04,
 -0.885942102175E-05,
 -0.447991560607E-05,
 -0.207963594384E-05,
 -0.111067675416E-05,
 -0.138435856935E-05,
 -0.812701410824E-06,
  0.485645147702E-05,
  0.125436950529E-04,
  0.205835723762E-04,
 -0.492842126415E-04,
 -0.608401625890E-04,
  0.466507176427E-04,
  0.353101147437E-04,
  0.524209145920E-06,
 -0.104804749854E-04,
 -0.552840858333E-04,
  0.444843447618E-04,
  0.209867336615E-03,
 -0.187407483015E-04,
 -0.162344956775E-03,
  0.682834838507E-06,
 -0.124209345053E-04,
 -0.938558508053E-05,
  0.778364490789E-04,
  0.196604060209E-04,
 -0.776129110912E-04,
  0.150857415008E-04,
 -0.218653562347E-05,
  0.492482383534E-05,
  0.656799937326E-04,
 -0.132777213959E-04,
 -0.257932067241E-03,
 -0.243965247780E-04,
  0.208378222643E-03
);
end;
