-- 17.02.2015
