package initial is

constant mm_1:real:=  0.288058870532E-08;
constant dm_1:real:=  0.706010261432E-04;
constant mm_2:real:=  0.653087233995E-08;
constant dm_2:real:=  0.245685234375E-03;
constant fi1_1:real:=  0.997970744648    ;
constant fi1_2:real:=  0.999999999731    ;
constant fi2_1:real:=  0.569280444689E-10;
constant fi2_2:real:=  0.996567701520    ;
constant fi3_1:real:= -0.803900764657    ;
constant fi3_2:real:=  0.953682688426    ;
constant el1_1:real:= -0.211089068271E-11;
constant el1_2:real:= -0.706066545973E-01;
constant el2_1:real:=   60748.3863376    ;
constant el2_2:real:=   103011.432553    ;

end;
