package ca23_dat_135 is

constant ca23_type135:integer:=1;
constant ca23_inve135:integer:=2;
signal ca23_ord135:real_vector(1 to 3):=( 6.0, 4.0, 2.0);
signal ca23_fak135:real_vector(1 to 4):=( 0.985831178093E-01, 0.214896594093, 4.92915589046,  4481.94303317);
constant ca23_anz135:integer:=       105;
signal ca23_data135:real_vector(1 to 105):=
(
  0.542306933822    ,
 -0.740386842324E-06,
  0.720568821477E-02,
  0.322049295306E-05,
  0.751730271837E-03,
 -0.240942008668E-05,
 -0.289635058843E-03,
 -0.263995134137    ,
 -0.368925030515E-06,
 -0.635444030127E-02,
  0.899365225491E-06,
 -0.526524808956E-03,
 -0.584595263498E-06,
  0.150831817484E-03,
  0.110604501845    ,
  0.603462236089E-05,
  0.304515033060E-02,
 -0.210651777072E-04,
  0.207972242616E-02,
  0.152142520666E-04,
 -0.100321596850E-02,
 -0.452052745975E-01,
  0.279215414060E-06,
 -0.203439389771E-02,
 -0.618977517276E-06,
 -0.318804969001E-03,
  0.426464804814E-06,
  0.144029153398E-03,
  0.142602144522E-01,
 -0.505978107854E-05,
  0.146106460573E-02,
  0.173056561416E-04,
 -0.150090775054E-02,
 -0.124855058955E-04,
  0.776553486190E-03,
  0.143653423042E-02,
  0.743263436233E-08,
  0.160044959285E-04,
 -0.803228499034E-08,
  0.136308414496E-05,
  0.358475269886E-08,
 -0.416685385735E-06,
 -0.869240962651E-03,
  0.149896486146E-07,
  0.210511687194E-04,
 -0.131463793645E-06,
 -0.132389255812E-03,
  0.163761782358E-06,
  0.137461505640E-03,
  0.225311815912E-03,
 -0.102808220284E-07,
 -0.473868752980E-04,
  0.719913234608E-07,
  0.144560785278E-03,
 -0.943223743738E-07,
 -0.133544308105E-03,
  0.160414276689E-03,
 -0.213217950350E-07,
 -0.557561700802E-05,
  0.142686711065E-06,
  0.126730249496E-03,
 -0.172882345242E-06,
 -0.133819126760E-03,
 -0.148668789733E-03,
  0.920599679777E-08,
  0.237455209961E-04,
 -0.707459957331E-07,
 -0.137997942915E-03,
  0.947343264883E-07,
  0.129107675393E-03,
 -0.118399980562E-05,
  0.148987863962E-05,
 -0.222691783012E-06,
 -0.476777613627E-05,
 -0.738545457443E-07,
  0.331893366571E-05,
  0.449827968438E-07,
  0.862812226397E-05,
  0.805519865032E-08,
  0.120952198188E-04,
 -0.430996241931E-07,
 -0.527685857835E-04,
  0.519859641738E-07,
  0.563497499202E-04,
 -0.100520108361E-04,
 -0.747287930498E-05,
 -0.562686656129E-04,
  0.240410713435E-04,
  0.254202088471E-03,
 -0.168735569076E-04,
 -0.270868997931E-03,
  0.124514522026E-04,
 -0.849562699570E-08,
 -0.106374067860E-04,
  0.450571130951E-07,
  0.524567362206E-04,
 -0.542134889736E-07,
 -0.560572546756E-04,
 -0.778143380199E-05,
  0.598330282174E-05,
  0.550617735205E-04,
 -0.192727574471E-04,
 -0.253850925105E-03,
  0.135530454458E-04,
  0.270538608615E-03
);
end;
