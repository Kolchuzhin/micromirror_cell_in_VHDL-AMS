package ca13_dat_135 is

constant ca13_type135:integer:=1;
constant ca13_inve135:integer:=2;
signal ca13_ord135:real_vector(1 to 3):=( 6.0, 4.0, 2.0);
signal ca13_fak135:real_vector(1 to 4):=( 0.985831178093E-01, 0.214896594093, 4.92915589046,  25.8982724106);
constant ca13_anz135:integer:=       105;
signal ca13_data135:real_vector(1 to 105):=
(
  0.712787356737    ,
  0.181329103793    ,
 -0.198113083053E-01,
  0.415892797113E-02,
 -0.151607352349E-02,
  0.510117685739E-03,
 -0.864166175900E-04,
  0.131868405193    ,
 -0.964863444974E-02,
  0.398115891210E-02,
 -0.161012595883E-02,
 -0.155831400923E-03,
 -0.505275369194E-03,
  0.763004730461E-03,
 -0.308005577990E-02,
  0.909312617619E-03,
 -0.870699594639E-03,
  0.190077627663E-03,
  0.252001828837E-03,
  0.483567931544E-03,
 -0.493523236677E-03,
  0.218171862281E-03,
 -0.667409977826E-04,
 -0.124685131761E-03,
  0.240911943103E-04,
  0.667608381442E-03,
 -0.461344511120E-03,
 -0.607432879339E-04,
 -0.215073903340E-04,
  0.427256401124E-04,
 -0.461361171262E-04,
 -0.227514577258E-03,
  0.202995007468E-03,
  0.421073453121E-03,
 -0.407527390907E-03,
  0.421043739170E-03,
 -0.152582546212E-03,
  0.295524933266E-04,
 -0.116907881666E-04,
  0.762110224378E-05,
 -0.530978591088E-05,
  0.171817175012E-05,
  0.450020366778E-04,
 -0.319188189261E-04,
  0.275007409332E-04,
  0.197672245698E-04,
 -0.736138956303E-04,
 -0.616556252274E-05,
  0.457246664647E-04,
 -0.274712583003E-04,
  0.257605796649E-04,
 -0.454028101855E-04,
 -0.475117590783E-04,
  0.134975493679E-03,
  0.290002963160E-04,
 -0.866826479489E-04,
  0.791356979132E-05,
 -0.348437202025E-06,
 -0.184306680704E-04,
 -0.293786717880E-04,
  0.925340289760E-04,
  0.290117402543E-06,
 -0.513456418971E-04,
 -0.256017894342E-05,
 -0.949046209333E-05,
  0.386573585059E-04,
  0.587289537342E-04,
 -0.153324274249E-03,
 -0.230173708129E-04,
  0.885236170079E-04,
 -0.219671321382E-04,
  0.888337536338E-05,
 -0.456143959107E-05,
  0.199953090426E-05,
 -0.975055781182E-06,
  0.144042664115E-05,
 -0.881146608730E-06,
  0.501199192251E-05,
 -0.128719199357E-04,
  0.152322292782E-04,
  0.511509165282E-04,
 -0.358553110466E-04,
 -0.475130447340E-04,
  0.666396203235E-05,
  0.316745177112E-06,
  0.547183276670E-05,
 -0.502409854721E-04,
 -0.919932790212E-05,
  0.187353002643E-03,
 -0.278804373605E-04,
 -0.136419069101E-03,
  0.557359955382E-06,
  0.210499747075E-04,
 -0.504401682096E-05,
 -0.137018544679E-03,
 -0.179920498034E-05,
  0.147802958781E-03,
  0.451739993974E-04,
 -0.258999776157E-05,
 -0.395721259818E-07,
  0.810245745013E-04,
 -0.223151505586E-04,
 -0.327361592376E-03,
  0.754402584337E-04,
  0.275149243680E-03
);
end;
